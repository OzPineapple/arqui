../5/adder4bit/fulladder.vhdl