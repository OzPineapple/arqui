library ieee;
use ieee.std_logic.all;

entity rom is
	port();
end rom;
