../5/adder4bit/halfadder.vhdl