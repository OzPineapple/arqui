../5/adder4bit/logicxor.vhdl