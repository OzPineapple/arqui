library ieee;
use ieee.std_logic_1164;

entity ram is
	port(
		clock:		in		std_logic;
		reset:		in		std_logic;
		mode:		in		std_logic;
	);
end ram;

architecture arch of ram is
begin
		
end arch;
