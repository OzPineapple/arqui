../5/adder4bit/logicxnor.vhdl