../5/adder4bit/logicor.vhdl