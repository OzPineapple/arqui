../5/adder4bit/logicand.vhdl