util/test-mult8bit.vhdl