library iee;
use ieee.std_logic_1164.all;

package packageadder4bit00 is
	component xora
	end component;
	component fa00
	end component;
	component anda0
	end component;
	component xnora
	end component;
end packageadder4bit00;
