library ieee;
use ieee.std_logic_1164.all;

entity adder4bit is
	port(
		sel:	in std_logic;
		anum:	in	std_logic_vector(3 downto 0);
		bnum:	in	std_logic_vector(3 downto 0);
		led:	out std_logic;
		sum:	out	std_logic_vector(3 downto 0)
	);
end adder4bit;

architecture adder4bit_arch of adder4bit is
	component fulladder  is
		port(
			anum:	in	std_logic;
			bnum:	in	std_logic;
			cin:	in	std_logic;
			sum:	out	std_logic;
			cout:	out	std_logic
		);
	end component;
	component logicxor  is
		port(
			a:	in	std_logic;
			b:	in	std_logic;
			o:	out	std_logic
		);
	end component;
	component logicxnor is
		port(
			a:	in	std_logic;
			b:	in	std_logic;
			o:	out	std_logic
		);
	end component;
	component logicand  is
		port(
			a:	in	std_logic;
			b:	in	std_logic;
			o:	out	std_logic
		);
	end component;
	signal carry:	std_logic_vector(3 downto 0);
	signal bneg:	std_logic_vector(3 downto 0);
	signal sneg:	std_logic_vector(3 downto 0);
	signal cend:	std_logic;
begin
	rest0:	logicxor	port map( a => sel, b => bnum(0), o => bneg(0) );
	rest1:	logicxor	port map( a => sel, b => bnum(1), o => bneg(1) );
	rest2:	logicxor	port map( a => sel, b => bnum(2), o => bneg(2) );
	rest3:	logicxor	port map( a => sel, b => bnum(3), o => bneg(3) );
	sneg0:	fulladder	port map(anum => anum(0),	bnum => bneg(0),	cin => sel,			cout => carry(0),	sum => sneg(0) );
	sneg1:	fulladder	port map(anum => anum(1),	bnum => bneg(1),	cin => carry(0),	cout => carry(1),	sum => sneg(1) );
	sneg2:	fulladder	port map(anum => anum(2),	bnum => bneg(2),	cin => carry(1),	cout => carry(2),	sum => sneg(2) );
	sneg3:	fulladder	port map(anum => anum(3),	bnum => bneg(3),	cin => carry(2),	cout => carry(3),	sum => sneg(3) );
	ledh:	logicxor	port map( a => carry(3), b => carry(2), o => led  );
	idkw:	logicxnor	port map( a => carry(3), b => carry(2), o => cend );
	sum0:	logicand	port map( a => cend,	 b => sneg(0),	o => sum(0) );
	sum1:	logicand	port map( a => cend,	 b => sneg(1),	o => sum(1) );
	sum2:	logicand	port map( a => cend,	 b => sneg(2),	o => sum(2) );
	sum3:	logicand	port map( a => cend,	 b => sneg(3),	o => sum(3) );
end adder4bit_arch;
