library ieee;
use ieee.std_logic_1164.all;

entity countRead is
	port(
		);
end countRead;

architecture arch of countRead is
begin
	if( clock'event
end countRead;
